module Rsa256Wrapper (
        input         avm_rst,
        input         avm_clk,
        output  [4:0] avm_address,
        output        avm_read,
        input  [31:0] avm_readdata,
        output        avm_write,
        output [31:0] avm_writedata,
        input         avm_waitrequest
    );


endmodule
