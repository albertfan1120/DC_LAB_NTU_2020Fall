// rsa_qsys.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module rsa_qsys (
		input  wire  clk_clk,                        //                        clk.clk
		input  wire  reset_reset_n,                  //                      reset.reset_n
		input  wire  uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire  uart_0_external_connection_txd,  //                           .txd
		output wire [19:0] sram_addr,
		inout  wire [15:0] sram_data,
		output wire  sram_we_n,
		output wire  sram_ce_n,
		output wire  sram_oe_n,
		output wire  sram_lb_n,
		output wire  sram_ub_n,
		output wire [7:0] vga_r,
		output wire [7:0] vga_g,
		output wire [7:0] vga_b,
		output wire vga_blank_n,
		output wire vga_hs,
		output wire vga_vs,
		output wire vga_clk,
		output wire  [19:0] debug_wire,
		input  wire  [17:0] SW,
		input  wire CLK25_2,
		input  wire CLK75_6
	);

	wire         altpll_0_c0_clk;                           // altpll_0:c0 -> [mm_interconnect_0:altpll_0_c0_clk, rst_controller_001:clk, uart_0:clk, version1_0:avm_clk]
	wire  [31:0] version1_0_avalon_master_0_readdata;       // mm_interconnect_0:version1_0_avalon_master_0_readdata -> version1_0:avm_readdata
	wire         version1_0_avalon_master_0_waitrequest;    // mm_interconnect_0:version1_0_avalon_master_0_waitrequest -> version1_0:avm_waitrequest
	wire   [4:0] version1_0_avalon_master_0_address;        // version1_0:avm_address -> mm_interconnect_0:version1_0_avalon_master_0_address
	wire         version1_0_avalon_master_0_read;           // version1_0:avm_read -> mm_interconnect_0:version1_0_avalon_master_0_read
	wire         version1_0_avalon_master_0_write;          // version1_0:avm_write -> mm_interconnect_0:version1_0_avalon_master_0_write
	wire  [31:0] version1_0_avalon_master_0_writedata;      // version1_0:avm_writedata -> mm_interconnect_0:version1_0_avalon_master_0_writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;    // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;      // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;       // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;          // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer; // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;         // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;     // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> altpll_0:reset
	wire         rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> [mm_interconnect_0:version1_0_reset_sink_reset_bridge_in_reset_reset, uart_0:reset_n, version1_0:avm_rst]
	assign vga_clk = altpll_0_c0_clk;
	rsa_qsys_altpll_0 altpll_0 (
		.clk       (clk_clk),                        //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                               //             pll_slave.read
		.write     (),                               //                      .write
		.address   (),                               //                      .address
		.readdata  (),                               //                      .readdata
		.writedata (),                               //                      .writedata
		.c0        (altpll_0_c0_clk),//25m                //                    c0.clk
		.c1        (altpll_0_c1_clk),//75m                //                    c1.clk
		.c2        (altpll_0_c2_clk),//0.01M                //                    c2.clk
		.areset    (),                               //        areset_conduit.export
		.locked    (),                               //        locked_conduit.export
		.phasedone ()                                //     phasedone_conduit.export
	);

	rsa_qsys_uart_0 uart_0 (
		.clk           (altpll_0_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           ()                                           //                 irq.irq
	);

	Top version1_0 (
		.avm_address     (version1_0_avalon_master_0_address),     // avalon_master_0.address
		.avm_read        (version1_0_avalon_master_0_read),        //                .read
		.avm_readdata    (version1_0_avalon_master_0_readdata),    //                .readdata
		.avm_write       (version1_0_avalon_master_0_write),       //                .write
		.avm_writedata   (version1_0_avalon_master_0_writedata),   //                .writedata
		.avm_waitrequest (version1_0_avalon_master_0_waitrequest), //                .waitrequest
		.avm_clk         (altpll_0_c0_clk),                        //      clock_sink.clk
		.avm_rst         (rst_controller_001_reset_out_reset),      //      reset_sink.reset

		//
		.o_SRAM_ADDR(sram_addr),
	   .io_SRAM_DQ(sram_data),
		.o_SRAM_WE_N(sram_we_n),
		.o_SRAM_CE_N(sram_ce_n),
		.o_SRAM_OE_N(sram_oe_n),
		.o_SRAM_LB_N(sram_lb_n),
		.o_SRAM_UB_N(sram_ub_n),
		// VGA interface
		.VGA_R(vga_r),
		.VGA_G(vga_g),
		.VGA_B(vga_b),
		.VGA_BLANK_N(vga_blank_n),
		.VGA_HS(vga_hs),
		.VGA_VS(vga_vs),
		//
		.debug_wire(debug_wire),
		.vga_clk(vga_clk1),
		.CLK50(clk_clk),
		.pll_clk(altpll_1_c0_clk),
		.SW(SW),
		.CLK25_2(altpll_0_c0_clk),
		.CLK75_6(altpll_0_c1_clk),
		.CLK1M(altpll_0_c2_clk)
	);

	rsa_qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                   (altpll_0_c0_clk),                           //                                 altpll_0_c0.clk
		.version1_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),        // version1_0_reset_sink_reset_bridge_in_reset.reset
		.version1_0_avalon_master_0_address                (version1_0_avalon_master_0_address),        //                  version1_0_avalon_master_0.address
		.version1_0_avalon_master_0_waitrequest            (version1_0_avalon_master_0_waitrequest),    //                                            .waitrequest
		.version1_0_avalon_master_0_read                   (version1_0_avalon_master_0_read),           //                                            .read
		.version1_0_avalon_master_0_readdata               (version1_0_avalon_master_0_readdata),       //                                            .readdata
		.version1_0_avalon_master_0_write                  (version1_0_avalon_master_0_write),          //                                            .write
		.version1_0_avalon_master_0_writedata              (version1_0_avalon_master_0_writedata),      //                                            .writedata
		.uart_0_s1_address                                 (mm_interconnect_0_uart_0_s1_address),       //                                   uart_0_s1.address
		.uart_0_s1_write                                   (mm_interconnect_0_uart_0_s1_write),         //                                            .write
		.uart_0_s1_read                                    (mm_interconnect_0_uart_0_s1_read),          //                                            .read
		.uart_0_s1_readdata                                (mm_interconnect_0_uart_0_s1_readdata),      //                                            .readdata
		.uart_0_s1_writedata                               (mm_interconnect_0_uart_0_s1_writedata),     //                                            .writedata
		.uart_0_s1_begintransfer                           (mm_interconnect_0_uart_0_s1_begintransfer), //                                            .begintransfer
		.uart_0_s1_chipselect                              (mm_interconnect_0_uart_0_s1_chipselect)     //                                            .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
